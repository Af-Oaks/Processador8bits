module Soma1bitSai3(entrada,Saida);


input wire[2:0]entrada;
output wire[2:0]Saida;


assign Saida = entrada + 1;


endmodule
