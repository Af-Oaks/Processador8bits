module Soma2num(entrada1,entrada2,Saida);


input wire[7:0]entrada1,entrada2;
output wire[7:0]Saida;


assign Saida = entrada1 + entrada2;


endmodule

