module portaOr2(entrada1,entrada2,Saida);


input wire entrada1,entrada2;
output wire Saida;


assign Saida = entrada1 | entrada2 ;


endmodule

